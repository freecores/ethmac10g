/////////////////////////////////////////////////////////////////////////////
//
//		Name of module 
//              23/1/06 - So far Mentor Precision indicates the current system runs as 101 MHz.
//
/////////////////////////////////////////////////////////////////////////////
module TRANSMIT_TOP(
TX_DATA, 
TX_DATA_VALID, 
TX_CLK, 
RESET, 
TX_START, 
TX_ACK, 
TX_UNDERRUN, 
TX_IFG_DELAY,
RXTXLINKFAULT, 
LOCALLINKFAULT,
TXSTATREGPLUS,
TXD, 
TXC, 
FC_TRANS_PAUSEDATA, 
FC_TRANS_PAUSEVAL, 
FC_TX_PAUSEDATA,
FC_TX_PAUSEVALID,
TX_CFG_REG_VALUE,
TX_CFG_REG_VALID
);


/////////////////////////////////////////////////////////////////////////////
//
//		Input and output ports definitions
//
/////////////////////////////////////////////////////////////////////////////

//Input from user logic
input [63:0] TX_DATA;
input [7:0] TX_DATA_VALID; // To accept the data valid to be available
input TX_CLK;
input RESET;
input TX_START; // This signify the first frame of data
input TX_UNDERRUN; // this will cause an error to be injected into the data
input [7:0] TX_IFG_DELAY; // this will cause a delay in the ack signal

//input to transmit fault signals
input RXTXLINKFAULT;
input LOCALLINKFAULT;

input [31:0] TX_CFG_REG_VALUE;
input TX_CFG_REG_VALID;

//output to stat register
output [9:0] TXSTATREGPLUS; // a pulse for each reg for stats

//output to user logic
output TX_ACK; //Generated by a counter

//output to XGMII
output [63:0] TXD;
output [7:0] TXC;

//output [15:0] BYTE_COUNTER_OUT;

//Pause inputs
//Transmit pause frames
input [15:0] FC_TRANS_PAUSEDATA; //pause frame data
input FC_TRANS_PAUSEVAL; //pulse signal to indicate a pause frame to be sent

//apply pause timing
input [15:0] FC_TX_PAUSEDATA;
input FC_TX_PAUSEVALID;



/////////////////////////////////////////////////////////////////////////////
//
//		Definitions and parameters
//
/////////////////////////////////////////////////////////////////////////////

//possibility to put this in a package.

//opcode definitions
parameter PAUSE_OPCODE = 16'b1000100000001000; //8808
parameter  VLAN_OPCODE = 16'b1000000100000000; //8100

//frame size definitions
parameter VLAN_FRAME_SIZE = 16'b0000010111110010;//1522 bytes
parameter JUMBO_FRAME_SIZE = 16'b0010001100101000;//9000 bytes
parameter NORMAL_FRAME_SIZE = 16'b0000010111101110;//1518 bytes
parameter MIN_FRAME_SIZE = 16'b0000000000111100; //60 bytes


//Frame definition
parameter IDLE_FRAME = 8'b00000111; //only six preambles as the first preamble is converted into a start flag
parameter IDLE_FRAME_8BYTES = 64'b0000011100000111000001110000011100000111000001110000011100000111;
parameter START_SEQ = 64'b1010101110101010101010101010101010101010101010101010101011111011;
parameter LOCAL_FAULT_SEQ = 64'b0000000100000000000000000000000000000001000000000000000000000000;
parameter REMOTE_FAULT_SEQ = 64'b0000001000000000000000000000000000000010000000000000000000000000;
parameter START_FRAME = 8'b11111011; //only valid in frame 0
parameter TERMINATE_FRAME = 8'b11111101;
parameter SFD_FRAME = 8'b10101011;
parameter PREAMBLE_FRAME = 8'b10101010;
parameter ERROR_FRAME = 8'b11111110;


parameter SOURCE_ADDR = 48'h010101010101;
parameter DEST_ADDR = 48'h101010101010;

parameter PAUSE_FRAME_LENGTH = 8'h02;

//need a parameter for min frame gap.

//Link fault signalling
// send lane 0


/////////////////////////////////////////////////////////////////////////////
//
//		Registers and wires
//
/////////////////////////////////////////////////////////////////////////////


reg [15:0] length_register;
wire [15:0] BYTE_COUNTER;
reg PARALLEL_CNT;

wire [31:0] CRC_32_64;
wire [31:0] CRC_OUT;

reg [31:0] CRC_OUT_REG;

reg error_flag_int;
reg insert_error;
reg [63:0] tx_data_int;

reg [63:0] TXD;
reg [7:0] TXC;
reg start_CRC8;

reg [7:0] TX_DATA_VALID_REG;
reg [63:0] TX_DATA_REG;


reg [15:0] DELAY_ACK;

wire  TX_ACK;

reg FRAME_START;

reg [63:0] TXD_DEL1;
reg [63:0] TXD_DEL2;
reg [63:0] TXD_DEL3;
reg [63:0] TXD_DEL4;
reg [63:0] TXD_DEL5;
reg [63:0] TXD_DEL6;
reg [63:0] TXD_DEL7;
reg [63:0] TXD_DEL8;
reg [63:0] TXD_DEL9;
reg [63:0] TXD_DEL10;
reg [63:0] TXD_DEL11;
reg [63:0] TXD_DEL12;

reg [7:0] TXC_DEL1;
reg [7:0] TXC_DEL2;
reg [7:0] TXC_DEL3;
reg [7:0] TXC_DEL4;
reg [7:0] TXC_DEL5;
reg [7:0] TXC_DEL6;
reg [7:0] TXC_DEL7;
reg [7:0] TXC_DEL8;
reg [7:0] TXC_DEL9;
reg [7:0] TXC_DEL10;
reg [7:0] TXC_DEL11;
reg [7:0] TXC_DEL12;

reg [7:0] OVERFLOW_VALID;
reg [63:0] OVERFLOW_DATA; 


reg [63:0] TXD_PAUSE_DEL0;
reg [63:0] TXD_PAUSE_DEL1;
reg [63:0] TXD_PAUSE_DEL2;
reg [63:0] TXD_PAUSE_DEL3;
reg [63:0] TXD_PAUSE_DEL4;
reg [63:0] TXD_PAUSE_DEL5;
reg [63:0] TXD_PAUSE_DEL6;
reg [63:0] TXD_PAUSE_DEL7;
reg [63:0] TXD_PAUSE_DEL8;

reg [7:0] TXC_PAUSE_DEL0;
reg [7:0] TXC_PAUSE_DEL1;
reg [7:0] TXC_PAUSE_DEL2;
reg [7:0] TXC_PAUSE_DEL3;
reg [7:0] TXC_PAUSE_DEL4;
reg [7:0] TXC_PAUSE_DEL5;
reg [7:0] TXC_PAUSE_DEL6;
reg [7:0] TXC_PAUSE_DEL7;
reg [7:0] TXC_PAUSE_DEL8;

/////////////////////////////////////////////////////////////////////////////
//
//		Start of code
//
/////////////////////////////////////////////////////////////////////////////




//TODO

//RX side. need to be able to receive data and calculate the CRC switching between 64 and 8 bit datapath.
//Therefore, the data need to be counted correctly.
//ERROR checking module or process will be needed. This will check if frame is correct length.
//Need to be able to remove redundant frames or columns and also padding. The error module will
//also check the tx_underrun signal as well.

//need to be able to cut-off bytes. 

//Need to add the link fault signalling and config registers.


//TX side. need to be able to insert the CRC with the data.
//need to define the first column of txd which is START 6 PRE and SFD.
//need to be able invert data_valid for txc.
//need to be able to transmit IDLEs.


//Format of output
//IDLE 07, START FB TERMINATE FD SFD 10101011 PREAMBLE 10101010  ERROR FE.

//IDLE START PREAMBLE SFD DA SA L/T DATA TERMINATE IDLE





integer i;
reg FRAME_START_DEL;
reg START_CRC8_DEL;
reg LOAD_CRC;
wire load_CRC8;
reg load_CRC8_del;
reg [3:0] APPEND_CRC_COUNT;
reg [15:0] CRC8_COUNT;

reg LOAD_OVERFLOW;

reg start_CRC8_count;

reg apply_pause_delay;

reg [63:0] store_data;
reg [7:0] store_valid;
reg [31:0] store_CRC;
reg [31:0] store_byte_count;
reg [15:0] store_pause_frame;

reg APPLY_CRC_SET;

reg [15:0] MAX_FRAME_SIZE;

reg [15:0] DATA_SIZE;


reg transmit_pause_frame;
reg PAUSEVAL_DEL;
reg PAUSEVAL_DEL1;
reg PAUSEVAL_DEL2;
wire RESET_ERR_PAUSE;
reg [15:0] store_transmit_pause_value;
reg [3:0] pause_frame_counter;
reg [63:0] shift_pause_data;
reg [7:0] shift_pause_valid;
wire transmit_pause_frame_valid;
reg append_start_pause;
reg append_start_pause_del;
reg transmit_pause_frame_del;

/////////////////////////////////////////////////////////////////////////////
//
//		Ack counter
//
/////////////////////////////////////////////////////////////////////////////


//Ack counter. need to be able to load the frame length, pause frame inter frame delay into the ack counter
// as this will delay the ack signal. The ack signal will initiate the rest of the data transmission from the
// user logic.

//need to stop the ack signal from transmitting when a PAUSE frame is transmitting

// Connect DUT to test bench 
//This seem to be one of the culprit for the timing violation
ack_counter U_ACK_CNT(
.clock(TX_CLK),
.reset(RESET),	
.ready(FRAME_START |START_CRC8_DEL | start_CRC8 | transmit_pause_frame),
.tx_start(TX_START),
.max_count(DELAY_ACK),
.tx_ack(TX_ACK)
);


//CRC for 64 bit data
//This seem to be one of the culprit for the timing violation
CRC32_D64 U_CRC64(
.DATA_IN(TX_DATA_REG), //need to swap between pause data
.CLK(TX_CLK),	
.RESET(RESET | TX_ACK | append_start_pause),
.START(FRAME_START | transmit_pause_frame_valid),
.CRC_OUT(CRC_32_64) //need to switch to output some how for a pause frame
);


//CRC for 8 bit data
CRC32_D8 U_CRC8(
.DATA_IN(tx_data_int), //8bit data
.CLK(TX_CLK),
.RESET(RESET),
.START(start_CRC8),  //this signal will be use to start
.LOAD(load_CRC8), //use this to load first
.CRC_IN(CRC_32_64),
.CRC_OUT(CRC_OUT)
);



//The start signal need to be high for the count
//This seem to be one of the culprit for the timing violation
byte_count_module U_byte_count_module(
.CLK(TX_CLK),
.RESET(RESET | TX_ACK),
.START(FRAME_START),
.PARALLEL_CNT(PARALLEL_CNT), //May need to remove as I don't require it
.BYTE_COUNTER(BYTE_COUNTER)
);


/////////////////////////////////////////////////////////////////////////////
//
//Still need to add more config stuff here!!!!!! For configuration register
//
/////////////////////////////////////////////////////////////////////////////

//Need to modify this to be setup by the config register
always @(posedge TX_CLK or posedge RESET)
begin
  if (RESET) begin
    APPLY_CRC_SET <= 0;
  end

end

//Need to expand to be setup by the config register
always @(posedge TX_CLK or posedge RESET)
begin
  if (RESET) begin
    MAX_FRAME_SIZE <= 1514;
  end
end

//Need to modify this to look for length in VLAN frame.
always @(posedge TX_CLK or posedge RESET)
begin
   if (RESET) begin
      length_register <= 0;
   end
   else if (BYTE_COUNTER == 8) begin
      length_register <= TX_DATA_REG[47:32];
   end
end
/////////////////////////////////////////////////////////////////////////////


/////////////////////////////////////////////////////////////////////////////
//
//	PAUSE FRAME
//
/////////////////////////////////////////////////////////////////////////////

always @(posedge TX_CLK)
begin
  PAUSEVAL_DEL <= FC_TRANS_PAUSEVAL;
  PAUSEVAL_DEL1 <= PAUSEVAL_DEL;
  PAUSEVAL_DEL2 <= PAUSEVAL_DEL1;
end

always @(posedge TX_CLK or posedge RESET)
begin
  if (RESET) begin
    transmit_pause_frame <= 0;
  end
  else if (PAUSEVAL_DEL2) begin
    transmit_pause_frame <= 1;
  end 
  else if (pause_frame_counter == 8) begin
    transmit_pause_frame <= 0;
  end 
end

always @(posedge TX_CLK or posedge RESET)
begin
  if (RESET) begin
    TXD_PAUSE_DEL0 <= 0;
    TXD_PAUSE_DEL1 <= 0;
    TXD_PAUSE_DEL2 <= 0;
    TXD_PAUSE_DEL3 <= 0;
    TXD_PAUSE_DEL4 <= 0;
    TXD_PAUSE_DEL5 <= 0;
    TXD_PAUSE_DEL6 <= 0;
    TXD_PAUSE_DEL7 <= 0;
    TXD_PAUSE_DEL8 <= 0;

    TXC_PAUSE_DEL0 <= 0;
    TXC_PAUSE_DEL1 <= 0;
    TXC_PAUSE_DEL2 <= 0;
    TXC_PAUSE_DEL3 <= 0;
    TXC_PAUSE_DEL4 <= 0; 
    TXC_PAUSE_DEL5 <= 0;
    TXC_PAUSE_DEL6 <= 0;
    TXC_PAUSE_DEL7 <= 0;
    TXC_PAUSE_DEL8 <= 0;

    store_transmit_pause_value <= 0;
  end
  else if (FC_TRANS_PAUSEVAL) begin
    store_transmit_pause_value <= FC_TRANS_PAUSEDATA;
    TXD_PAUSE_DEL1 <= {DEST_ADDR, SOURCE_ADDR[47:32]};
    TXD_PAUSE_DEL2 <= {SOURCE_ADDR[31:0], PAUSE_FRAME_LENGTH, PAUSE_OPCODE, FC_TRANS_PAUSEDATA};

    TXC_PAUSE_DEL1 <= 8'hff;
    TXC_PAUSE_DEL2 <= 8'hff;
    TXC_PAUSE_DEL3 <= 8'hff;
    TXC_PAUSE_DEL4 <= 8'hff; 
    TXC_PAUSE_DEL5 <= 8'hff;
    TXC_PAUSE_DEL6 <= 8'hff;
    TXC_PAUSE_DEL7 <= 8'hff;
    TXC_PAUSE_DEL8 <= 8'h0f;
  end 
end


always @(posedge TX_CLK or posedge RESET)
begin
  if (RESET) begin
    pause_frame_counter <= 0;
  end
  else if (transmit_pause_frame & !FRAME_START) begin
    pause_frame_counter <= pause_frame_counter + 1;
  end 
end


always @(posedge TX_CLK or posedge RESET)
begin
  if (RESET) begin
    shift_pause_data <= 0;
    shift_pause_valid <= 0;
  end
  else if (transmit_pause_frame & !FRAME_START) begin
    if (pause_frame_counter == 0) begin
      shift_pause_data <= TXD_PAUSE_DEL1;
    end
    else if (pause_frame_counter == 1) begin
      shift_pause_data <= TXD_PAUSE_DEL2;
    end
    else begin
      shift_pause_data <= 0;
    end 
    
    
    if (pause_frame_counter == 7) begin
      shift_pause_valid <= 8'h0f;
    end
    else if (pause_frame_counter < 7) begin
      shift_pause_valid <= 8'hff;
    end
    else begin
      shift_pause_valid <= 0;
    end 
  end
  else begin
    shift_pause_data <= 0;
    shift_pause_valid <= 0;
  end 
end





/////////////////////////////////////////////////////////////////////////////




//Signal that data is being processed and finshed.
always @(RESET or TX_ACK or TX_DATA_VALID_REG)
begin
  if (RESET) begin
     FRAME_START <= 0;
  end
  else if (TX_ACK) begin
     FRAME_START <= 1;
  end
  else if (TX_DATA_VALID_REG != 8'hff) begin
     FRAME_START <= 0;
  end
end


//Load the delay value for the acknowledge signal
always @(posedge TX_CLK or posedge RESET)
begin
   if (RESET) begin
     DELAY_ACK <= 16'h0001;
   end
   else if (apply_pause_delay) begin
     DELAY_ACK <= store_pause_frame;
   end
 end

//use for delaying the ack signal when pause is required
always @(posedge TX_CLK or posedge RESET)
begin
   if (RESET | TX_ACK) begin
     apply_pause_delay <= 0;
     store_pause_frame <= 0;
   end
   else if (FC_TX_PAUSEVALID) begin
     apply_pause_delay <= 1;
     store_pause_frame <= FC_TX_PAUSEDATA;
   end
end

//Shift valid into the system and also ensuring min frame is achieved
always @(posedge TX_CLK or posedge RESET)
begin
  if (RESET) begin
   
   TX_DATA_VALID_REG <= 0;
  end
  else if (FRAME_START) begin
   if (BYTE_COUNTER < 56) begin
     TX_DATA_VALID_REG <= 8'b11111111;
   end
   else if (BYTE_COUNTER == 56) begin
     TX_DATA_VALID_REG <= 8'b00001111 | TX_DATA_VALID;
   end
   else begin
     TX_DATA_VALID_REG <= TX_DATA_VALID;
   end
  end
  else if (transmit_pause_frame_valid) begin
     TX_DATA_VALID_REG <= shift_pause_valid;
  end
  else begin
   
   TX_DATA_VALID_REG <= 0;
  end

end


//Shifting data to the system. Also ensuring min frame is achieved
always @(posedge TX_CLK or posedge RESET)
begin
  if (RESET) begin
     TX_DATA_REG <= IDLE_FRAME_8BYTES;
  end
  else if (FRAME_START) begin
     if (BYTE_COUNTER < 56) begin
        case (TX_DATA_VALID)
      	8'b00000000 : begin
                      TX_DATA_REG <= 0;
                    end
        8'b00000001 : begin
                      TX_DATA_REG <= {56'h00000000000000, TX_DATA[7:0]};
                    end
        8'b00000011 : begin
                      TX_DATA_REG <= {48'h000000000000, TX_DATA[15:0]};
                    end                                                   
      	8'b00000111 : begin
                      TX_DATA_REG <= {40'h0000000000, TX_DATA[23:0]};
                    end
        8'b00001111 : begin
                      TX_DATA_REG <= {32'h00000000, TX_DATA[31:0]};
                    end
        8'b00011111 : begin
                      TX_DATA_REG <= {24'h000000, TX_DATA[39:0]};
                    end    
      	8'b00111111 : begin
                      TX_DATA_REG <= {16'h0000, TX_DATA[47:0]};
                    end
        8'b01111111 : begin
                      TX_DATA_REG <= {8'h00, TX_DATA[55:0]};
                    end
        8'b11111111 : begin
                      TX_DATA_REG <= TX_DATA;
                    end                    
        endcase                          
     end
     else if (BYTE_COUNTER == 56) begin
        TX_DATA_REG <= 0;
     end
     else begin
        TX_DATA_REG <= TX_DATA;
     end
  end
  else if (transmit_pause_frame_valid) begin
     TX_DATA_REG <= shift_pause_data;
  end  
  else begin
     TX_DATA_REG <= IDLE_FRAME_8BYTES;
  end

end



always @(posedge TX_CLK)
begin
   PARALLEL_CNT <= 1;
end


//Use for shifting data to CRC and loading start value for CRC
always @(posedge TX_CLK)
begin
  FRAME_START_DEL <= FRAME_START;
  transmit_pause_frame_del <= transmit_pause_frame;
  append_start_pause <= (!transmit_pause_frame_del & transmit_pause_frame);
  append_start_pause_del <= append_start_pause;
end

assign transmit_pause_frame_valid = (transmit_pause_frame_del & transmit_pause_frame);

assign RESET_ERR_PAUSE = (transmit_pause_frame_del & !transmit_pause_frame);
assign load_CRC8 = (FRAME_START_DEL & !FRAME_START) | (transmit_pause_frame_del & !transmit_pause_frame);





//store 64 bit data CRC result, data_valid, data
always @(posedge TX_CLK or posedge RESET)
begin
  if (RESET) begin
    store_data <= 0;
    store_valid <= 0;
    store_CRC <= 0;
    tx_data_int <= 0;
    store_byte_count <= 0;
  end
  else if (load_CRC8) begin
    store_data <= TX_DATA_REG;
    store_valid <= TX_DATA_VALID_REG;
    store_CRC <= CRC_32_64;
    store_byte_count <= BYTE_COUNTER;
  end
  else begin
    store_valid[6:0] <= store_valid[7:1];
    tx_data_int <= store_data[7:0];
    store_data[55:0] <= store_data[63:8];
  end
end





//Start CRC8 and load CRC8
always @(posedge TX_CLK or posedge RESET)
begin
  if (RESET) begin
    start_CRC8 <= 0;
    START_CRC8_DEL <= 0;
    error_flag_int <= 0;
  end
  else begin
    start_CRC8 <= store_valid[0];
    START_CRC8_DEL <= start_CRC8;
    if (load_CRC8 == 1 & TX_DATA_VALID_REG == 8'h00) begin
      error_flag_int  <= load_CRC8;
    end
    else begin
      error_flag_int <= START_CRC8_DEL & !start_CRC8;
    end
    
  end
end

//Use for determining the number of bytes in the data
always @(posedge TX_CLK or posedge RESET)
begin
  if (RESET) begin
     CRC8_COUNT <= 0;
  end
  else if (load_CRC8) begin
     CRC8_COUNT <= BYTE_COUNTER;
  end
  else if (start_CRC8) begin
     CRC8_COUNT <= CRC8_COUNT + 1;
  end
end

//Flag use for appending CRC and terminate
always @(APPEND_CRC_COUNT)
begin
  if (APPEND_CRC_COUNT == 9) begin
    LOAD_CRC <= 1;
  end
  else begin
    LOAD_CRC <= 0;
  end
end

//Flag use for appending CRC and terminate
always @(APPEND_CRC_COUNT)
begin
  if (APPEND_CRC_COUNT == 10) begin
    LOAD_OVERFLOW <= 1;
  end
  else begin
    LOAD_OVERFLOW <= 0;
  end
end

//Start the append counter
always @(posedge TX_CLK or posedge RESET)
begin
  if (RESET) begin
    start_CRC8_count <= 0;
  end
  else if (load_CRC8) begin
    start_CRC8_count <= 1;
  end
  else if (APPEND_CRC_COUNT == 10) begin
    start_CRC8_count <= 0;
  end
end

//Counter use to determine when to append CRC
always @(posedge TX_CLK or posedge RESET)
begin
  if (RESET | load_CRC8) begin
    APPEND_CRC_COUNT <= 0;
  end
  else if (start_CRC8_count) begin
    APPEND_CRC_COUNT <= APPEND_CRC_COUNT +1;
  end
end


//Append CRC and Terminate - still need to create non-crc version. Require a flag to stop CRC from generating.
always @(posedge TX_CLK or posedge RESET)
begin
  if (RESET) begin
    TXD_DEL1 <= 0;
    TXD_DEL2 <= 0;
    TXD_DEL3 <= 0; 
    TXD_DEL4 <= 0;
    TXD_DEL5 <= 0;
    TXD_DEL6 <= 0;
    TXD_DEL7 <= 0;
    TXD_DEL8 <= 0;
    TXD_DEL9 <= 0;
    TXD_DEL10 <= 0;
    TXD_DEL11 <= 0;
    TXD_DEL12 <= 0;
    TXC_DEL1 <= 0;
    TXC_DEL2 <= 0;
    TXC_DEL3 <= 0;
    TXC_DEL4 <= 0;
    TXC_DEL5 <= 0;
    TXC_DEL6 <= 0;
    TXC_DEL7 <= 0;
    TXC_DEL8 <= 0;
    TXC_DEL9 <= 0;
    TXC_DEL10 <= 0;
    TXC_DEL11 <= 0;     
    TXC_DEL12 <= 0; 
  end
  else begin
   
    //Append start seq.
    if (TX_ACK) begin
      TXD_DEL1 <= START_SEQ;
    end 
    else if (append_start_pause) begin
      TXD_DEL1 <= START_SEQ;
    end
    else begin
      TXD_DEL1 <= TX_DATA_REG;
    end
    
    TXD_DEL2 <= TXD_DEL1;
    TXD_DEL3 <= TXD_DEL2; 
    TXD_DEL4 <= TXD_DEL3;
    TXD_DEL5 <= TXD_DEL4;
    TXD_DEL6 <= TXD_DEL5;
    TXD_DEL7 <= TXD_DEL6;
    TXD_DEL8 <= TXD_DEL7;
    TXD_DEL9 <= TXD_DEL8;
    TXD_DEL10 <= TXD_DEL9;
    TXD_DEL11 <= TXD_DEL10;
    
    TXC_DEL1 <= TX_DATA_VALID_REG;
    TXC_DEL2 <= TXC_DEL1;
    TXC_DEL3 <= TXC_DEL2;
    TXC_DEL4 <= TXC_DEL3;
    TXC_DEL5 <= TXC_DEL4;
    TXC_DEL6 <= TXC_DEL5;
    TXC_DEL7 <= TXC_DEL6;
    TXC_DEL8 <= TXC_DEL7;
    TXC_DEL9 <= TXC_DEL8;
    TXC_DEL10 <= TXC_DEL9; 
    TXC_DEL11 <= TXC_DEL10;   
    
    if (LOAD_CRC) begin
    	case (TXC_DEL10)  
      	8'b00000000 : begin
                      TXD_DEL11[31:0] <= CRC_OUT[31:0];
                      if (insert_error) begin
                        TXD_DEL11[39:32] <= ERROR_FRAME;
                        TXD_DEL11[47:40] <= TERMINATE_FRAME;
                      end 
                      else begin
				TXD_DEL11[39:32] <= TERMINATE_FRAME;
                        TXD_DEL11[47:40] <= IDLE_FRAME;
                      end
                      
                      TXD_DEL11[55:48] <= IDLE_FRAME;
                      TXD_DEL11[63:56] <= IDLE_FRAME;
                      TXC_DEL11 <= 8'b00001111;
                      OVERFLOW_VALID <= 8'b00000000;
                      OVERFLOW_DATA <= IDLE_FRAME_8BYTES;                      
                    end
      	8'b00000001 : begin
		      TXD_DEL11[7:0] <= TXD_DEL10[7:0];
                      TXD_DEL11[39:8] <= CRC_OUT[31:0];
                      if (insert_error) begin
                        TXD_DEL11[47:40] <= ERROR_FRAME;
                        TXD_DEL11[55:48] <= TERMINATE_FRAME;
                      end 
                      else begin
                        TXD_DEL11[47:40] <= TERMINATE_FRAME;
                        TXD_DEL11[55:48] <= IDLE_FRAME;
                      end
                      TXD_DEL11[47:40] <= TERMINATE_FRAME;
                      TXD_DEL11[55:48] <= IDLE_FRAME;
                      TXD_DEL11[63:56] <= IDLE_FRAME;
                      TXD_DEL11 <= TXD_DEL10;
    		          TXC_DEL11 <= 8'b00011111;
                      OVERFLOW_VALID <= 8'b00000000;
                      OVERFLOW_DATA <= IDLE_FRAME_8BYTES;    		      
                    end
      	8'b00000011 : begin
		      TXD_DEL11[15:0] <= TXD_DEL10[15:0];
                      TXD_DEL11[47:16] <= CRC_OUT[31:0];
                      if (insert_error) begin
                        TXD_DEL11[55:48] <= ERROR_FRAME;
                        TXD_DEL11[63:56] <= TERMINATE_FRAME;
                      end 
                      else begin
                        TXD_DEL11[55:48] <= TERMINATE_FRAME;
                        TXD_DEL11[63:56] <= IDLE_FRAME;
                      end
                      TXC_DEL11 <= 8'b00111111;
                      OVERFLOW_VALID <= 8'b00000000;
                      OVERFLOW_DATA <= IDLE_FRAME_8BYTES; 	                
                    end
      	8'b00000111 : begin
		          TXD_DEL11[23:0] <= TXD_DEL10[23:0];
                      TXD_DEL11[55:24] <= CRC_OUT[31:0];
			    OVERFLOW_DATA <= IDLE_FRAME_8BYTES;
                      if (insert_error) begin
				TXD_DEL11[63:56] <= ERROR_FRAME;
				OVERFLOW_DATA[7:0] <= TERMINATE_FRAME;
                      end 
                      else begin
				TXD_DEL11[63:56] <= TERMINATE_FRAME;
                      end
                      TXC_DEL11 <= 8'b01111111;
                      OVERFLOW_VALID <= 8'b00000000;
                      OVERFLOW_DATA <= IDLE_FRAME_8BYTES;                      
                    end
      	8'b00001111 : begin
                      TXD_DEL11[31:0] <= TXD_DEL10[31:0];
		          TXD_DEL11[63:32]<= CRC_OUT[31:0];
	                TXC_DEL11<= 8'b11111111;
                      OVERFLOW_VALID <= 8'b00000000;
                      if (insert_error) begin
				OVERFLOW_DATA [7:0] <= ERROR_FRAME;
				OVERFLOW_DATA[15:8] <= TERMINATE_FRAME;
                      end 
                      else begin
				OVERFLOW_DATA [7:0]<= TERMINATE_FRAME; 
                        OVERFLOW_DATA [15:8]<= IDLE_FRAME; 
                      end
		      
                      OVERFLOW_DATA [23:16]<= IDLE_FRAME; 
                      OVERFLOW_DATA [31:24]<= IDLE_FRAME; 
                      OVERFLOW_DATA [39:32]<= IDLE_FRAME; 
                      OVERFLOW_DATA [47:40]<= IDLE_FRAME; 
                      OVERFLOW_DATA [55:48]<= IDLE_FRAME; 
                      OVERFLOW_DATA [63:56]<= IDLE_FRAME; 
                    end
      	8'b00011111 : begin
                      TXD_DEL11[39:0] <= TXD_DEL10[39:0];
                      TXD_DEL11[63:40] <= CRC_OUT[23:0];
                      TXC_DEL11 <= 8'b11111111;
                      OVERFLOW_VALID <= 8'b00000001;
		          OVERFLOW_DATA [7:0]<= CRC_OUT[31:24];
                      if (insert_error) begin
				OVERFLOW_DATA [15:8]<= ERROR_FRAME; 
                        OVERFLOW_DATA [23:16]<= TERMINATE_FRAME;
                      end 
                      else begin
				OVERFLOW_DATA [15:8]<= TERMINATE_FRAME; 
                        OVERFLOW_DATA [23:16]<= IDLE_FRAME;
                      end
                      OVERFLOW_DATA [31:24]<= IDLE_FRAME; 
                      OVERFLOW_DATA [39:32]<= IDLE_FRAME; 
                      OVERFLOW_DATA [47:40]<= IDLE_FRAME; 
                      OVERFLOW_DATA [55:48]<= IDLE_FRAME; 
                      OVERFLOW_DATA [63:56]<= IDLE_FRAME; 
                    end
      	8'b00111111 : begin
                      TXD_DEL11[47:0] <= TXD_DEL10[47:0];
                      TXD_DEL11[63:48] <= CRC_OUT[15:0];
                      TXC_DEL11 <= 8'b11111111;
                      OVERFLOW_VALID <= 8'b00000011;
		          OVERFLOW_DATA [15:0]<= CRC_OUT[31:16];  
                      if (insert_error) begin
				OVERFLOW_DATA [23:16]<= ERROR_FRAME; 
                        OVERFLOW_DATA [31:24]<= TERMINATE_FRAME;  
                      end 
                      else begin
				OVERFLOW_DATA [23:16]<= TERMINATE_FRAME; 
                        OVERFLOW_DATA [31:24]<= IDLE_FRAME; 
                      end                      
			    
                      OVERFLOW_DATA [39:32]<= IDLE_FRAME; 
                      OVERFLOW_DATA [47:40]<= IDLE_FRAME; 
                      OVERFLOW_DATA [55:48]<= IDLE_FRAME; 
                      OVERFLOW_DATA [63:56]<= IDLE_FRAME; 

                    end
      	8'b01111111 : begin
                      TXD_DEL11[55:0] <= TXD_DEL10[55:0];
                      TXD_DEL11[63:56] <= CRC_OUT[7:0];
                      TXC_DEL11 <= 8'b11111111;
                      OVERFLOW_VALID <= 8'b00000111;
		          OVERFLOW_DATA [23:0]<= CRC_OUT[31:8];  
                      if (insert_error) begin
				OVERFLOW_DATA [31:24]<= ERROR_FRAME; 
                        OVERFLOW_DATA [39:32]<= IDLE_FRAME;
                      end 
                      else begin
				OVERFLOW_DATA [31:24]<= TERMINATE_FRAME; 
                        OVERFLOW_DATA [39:32]<= IDLE_FRAME;
                      end
                       
                      OVERFLOW_DATA [47:40]<= IDLE_FRAME; 
                      OVERFLOW_DATA [55:48]<= IDLE_FRAME; 
                      OVERFLOW_DATA [63:56]<= IDLE_FRAME; 
                    end

      	endcase
    
    	
    
    end
    else if (LOAD_OVERFLOW) begin
	TXC_DEL11 <= OVERFLOW_VALID; 
        TXD_DEL11 <= OVERFLOW_DATA;    
    end
    
    
    TXD_DEL12 <= TXD_DEL11;
    TXC <= TXC_DEL12;
    TXD <= TXD_DEL12;    
    
  end
end



//Checking the data size from the byte count hence the -12 (remove address bytes)
always @(posedge TX_CLK or posedge RESET) 
begin
  if (RESET) begin
     DATA_SIZE <= 0;
  end
  else if (error_flag_int) begin
     DATA_SIZE <= CRC8_COUNT-12;
  end
end


//Indicate an error
always @(posedge TX_CLK or posedge RESET)
begin
  if (RESET | LOAD_OVERFLOW | RESET_ERR_PAUSE) begin
     insert_error <= 0;
  end
  else if (load_CRC8) begin
	if (length_register < MIN_FRAME_SIZE) begin
        if (CRC8_COUNT == 60) begin
     	    insert_error <= 0;
        end
        else begin
          insert_error <= 1;
        end
      end
      else if (length_register == DATA_SIZE) begin
	  if (CRC8_COUNT <= MAX_FRAME_SIZE) begin
     	    insert_error <= 0;
        end
        else begin
          insert_error <= 1;
        end
      end
      else begin
	  insert_error <= 1;
      end
  end
end


endmodule

